//OPT: -device TQFP44
//PIN: CHIP "top" ASSIGNED TO TQFP44
//PIN: O : 8
module top(output O);
  assign O = 1'b1;
endmodule
