module invert(input I, output O);
  INV n(.A(I), .QN(O));
endmodule
